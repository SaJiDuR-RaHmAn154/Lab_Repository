module subtractor (
    input wire [3:0] I,
    output wire [3:0] O
);
assign O = I - 1;    
endmodule


